`define WORD_LENGTH 32

